module kernel

pub fn kernel_main()
{
	
}